module ASR65(d_in, shamt, d_out); //module of Arthimetic Shift Right
	input	[64:0]	d_in; //input 
	input	[1:0]	shamt; 
	output [64:0] d_out; //output
	
	//instances 65 4to1 mux
	mx4 U0_mx4(d_in[0],d_in[1],d_in[2], d_in[3],shamt,d_out[0]);
	mx4 U1_mx4(d_in[1],d_in[2],d_in[3], d_in[4],shamt,d_out[1]);
	mx4 U2_mx4(d_in[2],d_in[3],d_in[4], d_in[5],shamt,d_out[2]);
	mx4 U3_mx4(d_in[3],d_in[4],d_in[5], d_in[6],shamt,d_out[3]);
	mx4 U4_mx4(d_in[4],d_in[5],d_in[6], d_in[7],shamt,d_out[4]);
	mx4 U5_mx4(d_in[5],d_in[6],d_in[7], d_in[8],shamt,d_out[5]);	
	mx4 U6_mx4(d_in[6],d_in[7],d_in[8], d_in[9],shamt,d_out[6]);
	mx4 U7_mx4(d_in[7],d_in[8],d_in[9], d_in[10],shamt,d_out[7]);
	mx4 U8_mx4(d_in[8],d_in[9],d_in[10], d_in[11],shamt,d_out[8]);
	mx4 U9_mx4(d_in[9],d_in[10],d_in[11], d_in[12],shamt,d_out[9]);
	mx4 U10_mx4(d_in[10],d_in[11],d_in[12], d_in[13],shamt,d_out[10]);
	mx4 U11_mx4(d_in[11],d_in[12],d_in[13], d_in[14],shamt,d_out[11]);
	mx4 U12_mx4(d_in[12],d_in[13],d_in[14], d_in[15],shamt,d_out[12]);
	mx4 U13_mx4(d_in[13],d_in[14],d_in[15], d_in[16],shamt,d_out[13]);	
	mx4 U14_mx4(d_in[14],d_in[15],d_in[16], d_in[17],shamt,d_out[14]);
	mx4 U15_mx4(d_in[15],d_in[16],d_in[17], d_in[18],shamt,d_out[15]);
	mx4 U16_mx4(d_in[16],d_in[17],d_in[18], d_in[19],shamt,d_out[16]);
	mx4 U17_mx4(d_in[17],d_in[18],d_in[19], d_in[20],shamt,d_out[17]);
	mx4 U18_mx4(d_in[18],d_in[19],d_in[20], d_in[21],shamt,d_out[18]);
	mx4 U19_mx4(d_in[19],d_in[20],d_in[21], d_in[22],shamt,d_out[19]);
	mx4 U20_mx4(d_in[20],d_in[21],d_in[22], d_in[23],shamt,d_out[20]);
	mx4 U21_mx4(d_in[21],d_in[22],d_in[23], d_in[24],shamt,d_out[21]);	
	mx4 U22_mx4(d_in[22],d_in[23],d_in[24], d_in[25],shamt,d_out[22]);
	mx4 U23_mx4(d_in[23],d_in[24],d_in[25], d_in[26],shamt,d_out[23]);
	mx4 U24_mx4(d_in[24],d_in[25],d_in[26], d_in[27],shamt,d_out[24]);
	mx4 U25_mx4(d_in[25],d_in[26],d_in[27], d_in[28],shamt,d_out[25]);
	mx4 U26_mx4(d_in[26],d_in[27],d_in[28], d_in[29],shamt,d_out[26]);
	mx4 U27_mx4(d_in[27],d_in[28],d_in[29], d_in[30],shamt,d_out[27]);
	mx4 U28_mx4(d_in[28],d_in[29],d_in[30], d_in[31],shamt,d_out[28]);
	mx4 U29_mx4(d_in[29],d_in[30],d_in[31], d_in[32],shamt,d_out[29]);	
	mx4 U30_mx4(d_in[30],d_in[31],d_in[32], d_in[33],shamt,d_out[30]);
	mx4 U31_mx4(d_in[31],d_in[32],d_in[33], d_in[34],shamt,d_out[31]);
	mx4 U32_mx4(d_in[32],d_in[33],d_in[34], d_in[35],shamt,d_out[32]);
	mx4 U33_mx4(d_in[33],d_in[34],d_in[35], d_in[36],shamt,d_out[33]);
	mx4 U34_mx4(d_in[34],d_in[35],d_in[36], d_in[37],shamt,d_out[34]);
	mx4 U35_mx4(d_in[35],d_in[36],d_in[37], d_in[38],shamt,d_out[35]);
	mx4 U36_mx4(d_in[36],d_in[37],d_in[38], d_in[39],shamt,d_out[36]);
	mx4 U37_mx4(d_in[37],d_in[38],d_in[39], d_in[40],shamt,d_out[37]);	
	mx4 U38_mx4(d_in[38],d_in[39],d_in[40], d_in[41],shamt,d_out[38]);
	mx4 U39_mx4(d_in[39],d_in[40],d_in[41], d_in[42],shamt,d_out[39]);
	mx4 U40_mx4(d_in[40],d_in[41],d_in[42], d_in[43],shamt,d_out[40]);
	mx4 U41_mx4(d_in[41],d_in[42],d_in[43], d_in[44],shamt,d_out[41]);
	mx4 U42_mx4(d_in[42],d_in[43],d_in[44], d_in[45],shamt,d_out[42]);
	mx4 U43_mx4(d_in[43],d_in[44],d_in[45], d_in[46],shamt,d_out[43]);
	mx4 U44_mx4(d_in[44],d_in[45],d_in[46], d_in[47],shamt,d_out[44]);
	mx4 U45_mx4(d_in[45],d_in[46],d_in[47], d_in[48],shamt,d_out[45]);	
	mx4 U46_mx4(d_in[46],d_in[47],d_in[48], d_in[49],shamt,d_out[46]);
	mx4 U47_mx4(d_in[47],d_in[48],d_in[49], d_in[50],shamt,d_out[47]);
	mx4 U48_mx4(d_in[48],d_in[49],d_in[50], d_in[51],shamt,d_out[48]);
	mx4 U49_mx4(d_in[49],d_in[50],d_in[51], d_in[52],shamt,d_out[49]);
	mx4 U50_mx4(d_in[50],d_in[51],d_in[52], d_in[53],shamt,d_out[50]);
	mx4 U51_mx4(d_in[51],d_in[52],d_in[53], d_in[54],shamt,d_out[51]);
	mx4 U52_mx4(d_in[52],d_in[53],d_in[54], d_in[55],shamt,d_out[52]);
	mx4 U53_mx4(d_in[53],d_in[54],d_in[55], d_in[56],shamt,d_out[53]);	
	mx4 U54_mx4(d_in[54],d_in[55],d_in[56], d_in[57],shamt,d_out[54]);
	mx4 U55_mx4(d_in[55],d_in[56],d_in[57], d_in[58],shamt,d_out[55]);
	mx4 U56_mx4(d_in[56],d_in[57],d_in[58], d_in[59],shamt,d_out[56]);
	mx4 U57_mx4(d_in[57],d_in[58],d_in[59], d_in[60],shamt,d_out[57]);
	mx4 U58_mx4(d_in[58],d_in[59],d_in[60], d_in[61],shamt,d_out[58]);
	mx4 U59_mx4(d_in[59],d_in[60],d_in[61], d_in[62],shamt,d_out[59]);
	mx4 U60_mx4(d_in[60],d_in[61],d_in[62], d_in[63],shamt,d_out[60]);
	mx4 U61_mx4(d_in[61],d_in[62],d_in[63], d_in[64],shamt,d_out[61]);	
	mx4 U62_mx4(d_in[62],d_in[63],d_in[64], d_in[64],shamt,d_out[62]);
	mx4 U63_mx4(d_in[63],d_in[64],d_in[64], d_in[64],shamt,d_out[63]);
	mx4 U64_mx4(d_in[64],d_in[64],d_in[64], d_in[64],shamt,d_out[64]);					
endmodule 