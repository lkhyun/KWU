module cla65(a,b,ci,s);
	input [64:0] a;
	input [64:0] b;
	input ci;
	output [64:0] s;
	wire [16:1] c;
	
cla4 U0_cla4(a[3:0],b[3:0],ci,c[1],s[3:0]);
cla4 U1_cla4(a[7:4],b[7:4],c[1],c[2],s[7:4]);
cla4 U2_cla4(a[11:8],b[11:8],c[2],c[3],s[11:8]);
cla4 U3_cla4(a[15:12],b[15:12],c[3],c[4],s[15:12]);
cla4 U4_cla4(a[19:16],b[19:16],c[4],c[5],s[19:16]);
cla4 U5_cla4(a[23:20],b[23:20],c[5],c[6],s[23:20]);
cla4 U6_cla4(a[27:24],b[27:24],c[6],c[7],s[27:24]);
cla4 U7_cla4(a[31:28],b[31:28],c[7],c[8],s[31:28]);
cla4 U8_cla4(a[35:32],b[35:32],c[8],c[9],s[35:32]);
cla4 U9_cla4(a[39:36],b[39:36],c[9],c[10],s[39:36]);
cla4 U10_cla4(a[43:40],b[43:40],c[10],c[11],s[43:40]);
cla4 U11_cla4(a[47:44],b[47:44],c[11],c[12],s[47:44]);
cla4 U12_cla4(a[51:48],b[51:48],c[12],c[13],s[51:48]);
cla4 U13_cla4(a[55:52],b[55:52],c[13],c[14],s[55:52]);
cla4 U14_cla4(a[59:56],b[59:56],c[14],c[15],s[59:56]);
cla4 U15_cla4(a[63:60],b[63:60],c[15],c[16],s[63:60]);
fa_v2 U16_fa_v2(a[64],b[64],c[16],s[64]); //1bit operate add

endmodule
